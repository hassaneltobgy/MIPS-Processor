--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:14:24 05/16/2022
-- Design Name:   
-- Module Name:   C:/Users/user/Desktop/Sophomore 2/Computer architecture/Major task/Ourcode/reg/Maincontroltb1.vhd
-- Project Name:  reg
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: controlunit
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Maincontroltb1 IS
END Maincontroltb1;
ARCHITECTURE behavior OF Maincontroltb1 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT controlunit
    PORT(
         opcode : IN  std_logic_vector(5 downto 0);
         output : OUT  std_logic_vector(10 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal opcode : std_logic_vector(5 downto 0) := (others => '0');

 	--Outputs
   signal output : std_logic_vector(10 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: controlunit PORT MAP (
          opcode => opcode,
          output => output
        );

   -- Clock process definitions
   <clock>_process :process
   begin
	<clock> <= '0';
	
	wait for <clock>_period/2;
	
	<clock> <= '1';
	wait for <clock>_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.      wait for 100 ns;	      wait for <clock>_period*10;
      -- insert stimulus here 

      wait;
   end process;

END;
