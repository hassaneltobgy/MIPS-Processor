
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use ieee.numeric_std.all;
entity Decoder is
    Port ( I : in  STD_LOGIC_VECTOR (4 downto 0);
			  E : in STD_LOGIC;
           O : out  STD_LOGIC_VECTOR (31 downto 0));
end Decoder;

architecture Behavioral of Decoder is

begin

O <= (OTHERS => 'Z') WHEN E = '0' ELSE

"00000000000000000000000000000001" WHEN I = "00000" ELSE --0
"00000000000000000000000000000010" WHEN I = "00001" ELSE --1
"00000000000000000000000000000100" WHEN I = "00010" ELSE --2
"00000000000000000000000000001000" WHEN I = "00011" ELSE  --3
"00000000000000000000000000010000" WHEN I = "00100" ELSE --4
"00000000000000000000000000100000" WHEN I = "00101" ELSE --5
"00000000000000000000000001000000" WHEN I = "00110" ELSE --6
"00000000000000000000000010000000" WHEN I = "00111" ELSE --7
"00000000000000000000000100000000" WHEN I = "01000" ELSE --8
"00000000000000000000001000000000" WHEN I = "01001" ELSE --9
"00000000000000000000010000000000" WHEN I = "01010" ELSE --10
"00000000000000000000100000000000" WHEN I = "01011" ELSE --11
"00000000000000000001000000000000" WHEN I = "01100" ELSE --12
"00000000000000000010000000000000" WHEN I = "01101" ELSE --13
"00000000000000000100000000000000" WHEN I = "01110" ELSE --14
"00000000000000001000000000000000" WHEN I = "01111" ELSE --15
"00000000000000010000000000000000" WHEN I = "10000" ELSE --16
"00000000000000100000000000000000" WHEN I = "10001" ELSE--17
"00000000000001000000000000000000" WHEN I = "10010" ELSE --18
"00000000000010000000000000000000" WHEN I = "10011" ELSE --19
"00000000000100000000000000000000" WHEN I = "10100" ELSE --20
"00000000001000000000000000000000" WHEN I = "10101" ELSE --21
"00000000010000000000000000000000" WHEN I = "10110" ELSE --22
"00000000100000000000000000000000" WHEN I = "10111" ELSE --23
"00000001000000000000000000000000" WHEN I = "11000" ELSE --24
"00000010000000000000000000000000" WHEN I = "11001" ELSE --25
"00000100000000000000000000000000" WHEN I = "11010" ELSE--26
"00001000000000000000000000000000" WHEN I = "11011" ELSE--27
"00010000000000000000000000000000" WHEN I = "11100" ELSE--28
"00100000000000000000000000000000" WHEN I = "11101" ELSE--29
"01000000000000000000000000000000" WHEN I = "11110" ELSE--30
"10000000000000000000000000000000" WHEN I = "11111" ELSE--31




(OTHERS => 'Z');
end behavioral;